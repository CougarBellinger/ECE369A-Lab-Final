`timescale 1ns / 1ps

module ForwardingUnit_tb();

reg Clk;
reg Reset;

wire 

endmodule